
module qsys (
	clk_clk,
	custom_logic_0_conduit_end_user_flag_1,
	custom_logic_0_conduit_end_user_flag_0,
	custom_logic_0_conduit_end_user_wrreq,
	custom_logic_0_conduit_end_user_data,
	custom_logic_0_conduit_end_user_wrclk);	

	input		clk_clk;
	output		custom_logic_0_conduit_end_user_flag_1;
	output		custom_logic_0_conduit_end_user_flag_0;
	input		custom_logic_0_conduit_end_user_wrreq;
	input	[31:0]	custom_logic_0_conduit_end_user_data;
	input		custom_logic_0_conduit_end_user_wrclk;
endmodule
